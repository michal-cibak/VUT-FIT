-- IVH Project: Patnáctka
-- Author: xcibak00 - Michal Cibák

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.std_logic_unsigned."conv_integer";


entity symbol_rom is
    port (
        ADDRESS : in std_logic_vector(3 downto 0);
        COLUMN  : in std_logic_vector(2 downto 0);
        ROW     : in std_logic_vector(2 downto 0);

        DATA    : out std_logic
    );
end symbol_rom;


architecture Behavioral of symbol_rom is
    type memory_t is array(0 to 15) of std_logic_vector(63 downto 0);
    constant MEMORY: memory_t := (
        (others => '0'),                                                    -- HOLE
        "0000000000111000000100000001000000010100000110000001000000000000", --  1
        "0000000000111100000001000001100000100000001001000001100000000000", --  2
        "0000000000011000001001000010000000010000001001000001100000000000", --  3
        "0000000000010000000100000011110000010100000001000000100000000000", --  4
        "0000000000011000001001000010000000011100000001000011110000000000", --  5
        "0000000000011000001001000010010000011100000001000011100000000000", --  6
        "0000000000001000000010000001000000010000001000000011110000000000", --  7
        "0000000000011000001001000010010000011000001001000001100000000000", --  8
        "0000000000011000001001000010000000111000001001000001100000000000", --  9
        "0000000000101110010101000101010001010100010101100010010000000000", -- 10
        "0000000001111110001001000010010000100100001101100010010000000000", -- 11
        "0000000001111110000101000010010001000100010101100010010000000000", -- 12
        "0000000000101110010101000100010000100100010001100011010000000000", -- 13
        "0000000000101110001001000111010000010100000101100010010000000000", -- 14
        "0000000000101110010101000100010000110100000101100111010000000000"  -- 15
    );

begin
    DATA <= MEMORY(conv_integer(ADDRESS))(conv_integer(ROW & COLUMN));
end Behavioral;
